library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity controlModule is 
  port (
    controlIn: in STD_LOGIC_VECTOR(31 downto 26);
    RegDst, Jump, Branch, MemRead, MemtoReg, MemWrite, ALUSrc, RegWrite: out STD_LOGIC;
    ALUOp: out STD_LOGIC_VECTOR(1 downto 0)
  );
end controlModule;
architecture behavioral of controlModule is
begin
control_process: process(controlIn)   
  begin
    if controlIn = "000000" then --add
      RegDst <= '1';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '1';
      ALUOp <= "10";
    elsif controlIn = "001000" then --addi
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00"; --uses lw/sw command ALUOp since this corresponds to add
    elsif controlIn = "001001" then --ALU needs modification to support unsigned addition
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "10";
    elsif controlIn = "001100" then --andi
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "10";
    elsif controlIn = "000100" then --beq
      RegDst <= '0';
      Jump <= '0';
      Branch <= '1';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "01";
    elsif controlIn = "000101" then --bne
      RegDst <= '0';
      Jump <= '0';
      Branch <= '1';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "11"; --assign unused ALUOp to this signal
    elsif controlIn = "000010" then --j
      RegDst <= '0';
      Jump <= '1';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "000011" then --jal
      RegDst <= '0';
      Jump <= '1';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "100100" then --lbu
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '1'; 
      MemtoReg <= '1'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "100101" then --lhu
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '1'; 
      MemtoReg <= '1'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "110000" then --ll
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '1'; 
      MemtoReg <= '1'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "001111" then --lui
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '1'; 
      MemtoReg <= '1'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "100011" then --lw
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '1'; 
      MemtoReg <= '1'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "001101" then --ori
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '1';
      ALUOp <= "00";
    elsif controlIn = "001010" then --slti
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "001011" then --sltiu
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "101000" then --sb
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '1'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "111000" then --sc
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '1'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "101001" then --sh
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '1'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    elsif controlIn = "101011" then --sw
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '1'; 
      ALUSrc <= '1'; 
      RegWrite <= '0';
      ALUOp <= "00";
    else
      RegDst <= '0';
      Jump <= '0';
      Branch <= '0';
      MemRead <= '0'; 
      MemtoReg <= '0'; 
      MemWrite <= '0'; 
      ALUSrc <= '0'; 
      RegWrite <= '0';
      ALUOp <= "00";
    end if; 
  end process control_process; 
end behavioral;    
